module Addcout4 (input [3:0] I0, input [3:0] I1, output [3:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
assign O = {inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst7_CO;
endmodule

module Register4 (input [3:0] I, output [3:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
assign O = {inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter4 (output [3:0] O, output  COUT, input  CLK);
wire [3:0] inst0_O;
wire  inst0_COUT;
wire [3:0] inst1_O;
Addcout4 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register4 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout3 (input [2:0] I0, input [2:0] I1, output [2:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
assign O = {inst4_O,inst2_O,inst0_O};
assign COUT = inst5_CO;
endmodule

module Register3CE (input [2:0] I, output [2:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
assign O = {inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter3CE (output [2:0] O, output  COUT, input  CLK, input  CE);
wire [2:0] inst0_O;
wire  inst0_COUT;
wire [2:0] inst1_O;
Addcout3 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register3CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout8 (input [7:0] I0, input [7:0] I1, output [7:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
assign O = {inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst15_CO;
endmodule

module Register8CE (input [7:0] I, output [7:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter8CE (output [7:0] O, output  COUT, input  CLK, input  CE);
wire [7:0] inst0_O;
wire  inst0_COUT;
wire [7:0] inst1_O;
Addcout8 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register8CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Invert8 (input [7:0] I, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst4 (.I0(I[4]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst5 (.I0(I[5]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst6 (.I0(I[6]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(I[7]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Register3CER (input [2:0] I, output [2:0] O, input  CLK, input  CE, input  RESET);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
SB_DFFESR inst0 (.C(CLK), .R(RESET), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFESR inst1 (.C(CLK), .R(RESET), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFESR inst2 (.C(CLK), .R(RESET), .E(CE), .D(I[2]), .Q(inst2_Q));
assign O = {inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter3CER (output [2:0] O, output  COUT, input  CLK, input  CE, input  RESET);
wire [2:0] inst0_O;
wire  inst0_COUT;
wire [2:0] inst1_O;
Addcout3 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register3CER inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE), .RESET(RESET));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module PISO8CE (input  SI, input [7:0] PI, input  LOAD, output  O, input  CLK, input  CE);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire [7:0] inst8_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(SI), .I1(PI[0]), .I2(LOAD), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(inst8_O[0]), .I1(PI[1]), .I2(LOAD), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(inst8_O[1]), .I1(PI[2]), .I2(LOAD), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(inst8_O[2]), .I1(PI[3]), .I2(LOAD), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(inst8_O[3]), .I1(PI[4]), .I2(LOAD), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(inst8_O[4]), .I1(PI[5]), .I2(LOAD), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(inst8_O[5]), .I1(PI[6]), .I2(LOAD), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(inst8_O[6]), .I1(PI[7]), .I2(LOAD), .I3(1'b0), .O(inst7_O));
Register8CE inst8 (.I({inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O}), .O(inst8_O), .CLK(CLK), .CE(CE));
assign O = inst8_O[7];
endmodule

module Addcout9 (input [8:0] I0, input [8:0] I1, output [8:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
wire  inst16_O;
wire  inst17_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst16 (.I0(1'b0), .I1(I0[8]), .I2(I1[8]), .I3(inst15_CO), .O(inst16_O));
SB_CARRY inst17 (.I0(I0[8]), .I1(I1[8]), .CI(inst15_CO), .CO(inst17_CO));
assign O = {inst16_O,inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst17_CO;
endmodule

module Register9CER (input [8:0] I, output [8:0] O, input  CLK, input  CE, input  RESET);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
SB_DFFESR inst0 (.C(CLK), .R(RESET), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFESR inst1 (.C(CLK), .R(RESET), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFESR inst2 (.C(CLK), .R(RESET), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFESR inst3 (.C(CLK), .R(RESET), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFESR inst4 (.C(CLK), .R(RESET), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFESR inst5 (.C(CLK), .R(RESET), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFESR inst6 (.C(CLK), .R(RESET), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFESR inst7 (.C(CLK), .R(RESET), .E(CE), .D(I[7]), .Q(inst7_Q));
SB_DFFESR inst8 (.C(CLK), .R(RESET), .E(CE), .D(I[8]), .Q(inst8_Q));
assign O = {inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter9CER (output [8:0] O, output  COUT, input  CLK, input  CE, input  RESET);
wire [8:0] inst0_O;
wire  inst0_COUT;
wire [8:0] inst1_O;
Addcout9 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register9CER inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE), .RESET(RESET));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Invert9 (input [8:0] I, output [8:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst4 (.I0(I[4]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst5 (.I0(I[5]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst6 (.I0(I[6]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(I[7]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst8 (.I0(I[8]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst8_O));
assign O = {inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Register8CER (input [7:0] I, output [7:0] O, input  CLK, input  CE, input  RESET);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFFESR inst0 (.C(CLK), .R(RESET), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFESR inst1 (.C(CLK), .R(RESET), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFESR inst2 (.C(CLK), .R(RESET), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFESR inst3 (.C(CLK), .R(RESET), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFESR inst4 (.C(CLK), .R(RESET), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFESR inst5 (.C(CLK), .R(RESET), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFESR inst6 (.C(CLK), .R(RESET), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFESR inst7 (.C(CLK), .R(RESET), .E(CE), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter8CER (output [7:0] O, output  COUT, input  CLK, input  CE, input  RESET);
wire [7:0] inst0_O;
wire  inst0_COUT;
wire [7:0] inst1_O;
Addcout8 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register8CER inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE), .RESET(RESET));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Invert4 (input [3:0] I, output [3:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
assign O = {inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Register4CER (input [3:0] I, output [3:0] O, input  CLK, input  CE, input  RESET);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
SB_DFFESR inst0 (.C(CLK), .R(RESET), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFESR inst1 (.C(CLK), .R(RESET), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFESR inst2 (.C(CLK), .R(RESET), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFESR inst3 (.C(CLK), .R(RESET), .E(CE), .D(I[3]), .Q(inst3_Q));
assign O = {inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter4CER (output [3:0] O, output  COUT, input  CLK, input  CE, input  RESET);
wire [3:0] inst0_O;
wire  inst0_COUT;
wire [3:0] inst1_O;
Addcout4 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register4CER inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE), .RESET(RESET));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module SIPO10CE (input  I, output [9:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(inst0_Q), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(inst1_Q), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(inst2_Q), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(inst3_Q), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(inst4_Q), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(inst5_Q), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(inst6_Q), .Q(inst7_Q));
SB_DFFE inst8 (.C(CLK), .E(CE), .D(inst7_Q), .Q(inst8_Q));
SB_DFFE inst9 (.C(CLK), .E(CE), .D(inst8_Q), .Q(inst9_Q));
assign O = {inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Mux2x4 (input [3:0] I0, input [3:0] I1, input  S, output [3:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(S), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(S), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(S), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(S), .I3(1'b0), .O(inst3_O));
assign O = {inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module main (output  D4, output  D5, output  D6, output  D7, input  O, output  I, output  D3, output  D2, output  D1, output  D0, input  CLKIN, input  RX);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire [3:0] inst3_O;
wire  inst3_COUT;
wire [2:0] inst4_O;
wire  inst4_COUT;
wire  inst5_O;
wire [7:0] inst6_O;
wire  inst6_COUT;
wire  inst7_O;
wire [7:0] inst8_O;
wire [7:0] inst9_O;
wire  inst9_COUT;
wire  inst10_Q;
wire [2:0] inst11_O;
wire  inst11_COUT;
wire  inst12_O;
wire  inst13_Q;
wire  inst14_O;
wire  inst15_O;
wire  inst16_O;
wire  inst17_O;
wire  inst18_O;
wire  inst19_O;
wire  inst20_O;
wire [8:0] inst21_O;
wire  inst21_COUT;
wire  inst22_O;
wire [8:0] inst23_O;
wire [8:0] inst24_O;
wire  inst24_COUT;
wire [8:0] inst25_O;
wire  inst25_COUT;
wire  inst26_Q;
wire  inst27_O;
wire  inst28_O;
wire [7:0] inst29_O;
wire  inst29_COUT;
wire  inst30_O;
wire  inst31_O;
wire  inst32_O;
wire  inst33_O;
wire  inst34_O;
wire  inst35_O;
wire  inst36_O;
wire  inst37_O;
wire  inst38_O;
wire  inst39_O;
wire  inst40_O;
wire  inst41_O;
wire  inst42_O;
wire  inst43_O;
wire  inst44_O;
wire  inst45_O;
wire  inst46_O;
wire  inst47_O;
wire  inst48_O;
wire  inst49_O;
wire  inst50_O;
wire  inst51_O;
wire  inst52_O;
wire  inst53_O;
wire  inst54_O;
wire  inst55_O;
wire  inst56_O;
wire  inst57_O;
wire  inst58_O;
wire  inst59_O;
wire  inst60_O;
wire  inst61_O;
wire  inst62_O;
wire  inst63_O;
wire  inst64_O;
wire  inst65_O;
wire  inst66_O;
wire  inst67_O;
wire  inst68_O;
wire  inst69_O;
wire  inst70_O;
wire  inst71_O;
wire  inst72_O;
wire  inst73_O;
wire  inst74_O;
wire  inst75_O;
wire  inst76_O;
wire  inst77_O;
wire  inst78_O;
wire  inst79_O;
wire  inst80_O;
wire  inst81_O;
wire  inst82_O;
wire  inst83_O;
wire  inst84_O;
wire  inst85_O;
wire  inst86_O;
wire  inst87_O;
wire  inst88_O;
wire  inst89_O;
wire  inst90_O;
wire  inst91_O;
wire  inst92_O;
wire  inst93_O;
wire  inst94_O;
wire  inst95_Q;
wire  inst96_O;
wire  inst97_O;
wire  inst98_O;
wire [3:0] inst99_O;
wire [3:0] inst100_O;
wire  inst100_COUT;
wire  inst101_O;
wire  inst102_O;
wire  inst103_O;
wire  inst104_O;
wire [3:0] inst105_O;
wire  inst105_COUT;
wire  inst106_O;
wire  inst107_O;
wire  inst108_O;
wire [9:0] inst109_O;
wire [15:0] inst110_RDATA;
wire [7:0] inst111_O;
wire  inst111_COUT;
wire  inst112_O;
wire  inst113_O;
wire  inst114_O;
wire  inst115_O;
wire  inst116_O;
wire  inst117_O;
wire  inst118_O;
wire  inst119_O;
wire  inst120_O;
wire  inst121_O;
wire  inst122_O;
wire  inst123_O;
wire  inst124_O;
wire  inst125_O;
wire  inst126_O;
wire  inst127_O;
wire  inst128_O;
wire  inst129_O;
wire  inst130_O;
wire  inst131_O;
wire  inst132_O;
wire  inst133_O;
wire  inst134_O;
wire  inst135_O;
wire  inst136_O;
wire  inst137_O;
wire  inst138_O;
wire  inst139_O;
wire  inst140_O;
wire  inst141_O;
wire  inst142_O;
wire  inst143_O;
wire  inst144_O;
wire [8:0] inst145_O;
wire  inst145_COUT;
wire [3:0] inst146_O;
wire  inst147_O;
wire [3:0] inst148_O;
wire [3:0] inst149_O;
wire  inst149_COUT;
wire  inst150_O;
SB_DFF inst0 (.C(CLKIN), .D(O), .Q(inst0_Q));
SB_DFF inst1 (.C(CLKIN), .D(inst0_Q), .Q(inst1_Q));
SB_DFF inst2 (.C(CLKIN), .D(inst1_Q), .Q(inst2_Q));
Counter4 inst3 (.O(inst3_O), .COUT(inst3_COUT), .CLK(CLKIN));
Counter3CE inst4 (.O(inst4_O), .COUT(inst4_COUT), .CLK(CLKIN), .CE(inst3_COUT));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst5 (.I0(inst3_COUT), .I1(inst4_COUT), .I2(1'b0), .I3(1'b0), .O(inst5_O));
Counter8CE inst6 (.O(inst6_O), .COUT(inst6_COUT), .CLK(CLKIN), .CE(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(inst9_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
Invert8 inst8 (.I({1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .O(inst8_O));
Addcout8 inst9 (.I0(inst6_O), .I1(inst8_O), .O(inst9_O), .COUT(inst9_COUT));
SB_DFFE inst10 (.C(CLKIN), .E(inst3_COUT), .D(inst7_O), .Q(inst10_Q));
Counter3CER inst11 (.O(inst11_O), .COUT(inst11_COUT), .CLK(CLKIN), .CE(inst3_COUT), .RESET(inst15_O));
SB_LUT4 #(.LUT_INIT(16'h0080)) inst12 (.I0(inst11_O[0]), .I1(inst11_O[1]), .I2(inst11_O[2]), .I3(1'b0), .O(inst12_O));
SB_DFFE inst13 (.C(CLKIN), .E(inst3_COUT), .D(inst14_O), .Q(inst13_Q));
SB_LUT4 #(.LUT_INIT(16'h5454)) inst14 (.I0(inst12_O), .I1(inst7_O), .I2(inst13_Q), .I3(1'b0), .O(inst14_O));
SB_LUT4 #(.LUT_INIT(16'h2222)) inst15 (.I0(inst12_O), .I1(inst13_Q), .I2(1'b0), .I3(1'b0), .O(inst15_O));
PISO8CE inst16 (.SI(1'b1), .PI({inst110_RDATA[0],inst110_RDATA[2],inst110_RDATA[4],inst110_RDATA[6],inst110_RDATA[8],inst110_RDATA[10],inst110_RDATA[12],inst110_RDATA[14]}), .LOAD(inst17_O), .O(inst16_O), .CLK(CLKIN), .CE(inst3_COUT));
SB_LUT4 #(.LUT_INIT(16'h2222)) inst17 (.I0(inst7_O), .I1(inst13_Q), .I2(1'b0), .I3(1'b0), .O(inst17_O));
SB_LUT4 #(.LUT_INIT(16'h4444)) inst18 (.I0(inst13_Q), .I1(inst3_COUT), .I2(1'b0), .I3(1'b0), .O(inst18_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst19 (.I0(inst13_Q), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst19_O));
SB_LUT4 #(.LUT_INIT(16'h8080)) inst20 (.I0(inst19_O), .I1(inst3_COUT), .I2(inst7_O), .I3(1'b0), .O(inst20_O));
Counter9CER inst21 (.O(inst21_O), .COUT(inst21_COUT), .CLK(CLKIN), .CE(inst20_O), .RESET(inst22_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst22 (.I0(inst24_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst22_O));
Invert9 inst23 (.I(inst21_O), .O(inst23_O));
Addcout9 inst24 (.I0({1'b0,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b1}), .I1(inst23_O), .O(inst24_O), .COUT(inst24_COUT));
Addcout9 inst25 (.I0(inst21_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst25_O), .COUT(inst25_COUT));
SB_DFF inst26 (.C(CLKIN), .D(inst2_Q), .Q(inst26_Q));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst27 (.I0(inst2_Q), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst27_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst28 (.I0(inst26_Q), .I1(inst27_O), .I2(1'b0), .I3(1'b0), .O(inst28_O));
Counter8CER inst29 (.O(inst29_O), .COUT(inst29_COUT), .CLK(CLKIN), .CE(1'b1), .RESET(inst62_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst30 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst30_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst31 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst31_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst32 (.I0(inst30_O), .I1(inst31_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst32_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst33 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst33_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst34 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst34_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst35 (.I0(inst33_O), .I1(inst34_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst35_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst36 (.I0(inst32_O), .I1(inst35_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst36_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst37 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst37_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst38 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst38_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst39 (.I0(inst37_O), .I1(inst38_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst39_O));
SB_LUT4 #(.LUT_INIT(16'h0040)) inst40 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst40_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst41 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst41_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst42 (.I0(inst40_O), .I1(inst41_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst42_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst43 (.I0(inst39_O), .I1(inst42_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst43_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst44 (.I0(inst36_O), .I1(inst43_O), .I2(inst29_O[6]), .I3(1'b0), .O(inst44_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst45 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst45_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst46 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst46_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst47 (.I0(inst45_O), .I1(inst46_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst47_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst48 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst48_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst49 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst49_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst50 (.I0(inst48_O), .I1(inst49_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst50_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst51 (.I0(inst47_O), .I1(inst50_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst51_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst52 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst52_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst53 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst53_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst54 (.I0(inst52_O), .I1(inst53_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst54_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst55 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst55_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst56 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst56_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst57 (.I0(inst55_O), .I1(inst56_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst57_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst58 (.I0(inst54_O), .I1(inst57_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst58_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst59 (.I0(inst51_O), .I1(inst58_O), .I2(inst29_O[6]), .I3(1'b0), .O(inst59_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst60 (.I0(inst44_O), .I1(inst59_O), .I2(inst29_O[7]), .I3(1'b0), .O(inst60_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst61 (.I0(inst60_O), .I1(inst28_O), .I2(1'b0), .I3(1'b0), .O(inst61_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst62 (.I0(inst61_O), .I1(1'b1), .I2(1'b0), .I3(1'b0), .O(inst62_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst63 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst63_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst64 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst64_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst65 (.I0(inst63_O), .I1(inst64_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst65_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst66 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst66_O));
SB_LUT4 #(.LUT_INIT(16'h0008)) inst67 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst67_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst68 (.I0(inst66_O), .I1(inst67_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst68_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst69 (.I0(inst65_O), .I1(inst68_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst69_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst70 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst70_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst71 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst71_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst72 (.I0(inst70_O), .I1(inst71_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst72_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst73 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst73_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst74 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst74_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst75 (.I0(inst73_O), .I1(inst74_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst75_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst76 (.I0(inst72_O), .I1(inst75_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst76_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst77 (.I0(inst69_O), .I1(inst76_O), .I2(inst29_O[6]), .I3(1'b0), .O(inst77_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst78 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst78_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst79 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst79_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst80 (.I0(inst78_O), .I1(inst79_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst80_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst81 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst81_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst82 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst82_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst83 (.I0(inst81_O), .I1(inst82_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst83_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst84 (.I0(inst80_O), .I1(inst83_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst84_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst85 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst85_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst86 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst86_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst87 (.I0(inst85_O), .I1(inst86_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst87_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst88 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst88_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst89 (.I0(inst29_O[0]), .I1(inst29_O[1]), .I2(inst29_O[2]), .I3(inst29_O[3]), .O(inst89_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst90 (.I0(inst88_O), .I1(inst89_O), .I2(inst29_O[4]), .I3(1'b0), .O(inst90_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst91 (.I0(inst87_O), .I1(inst90_O), .I2(inst29_O[5]), .I3(1'b0), .O(inst91_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst92 (.I0(inst84_O), .I1(inst91_O), .I2(inst29_O[6]), .I3(1'b0), .O(inst92_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst93 (.I0(inst77_O), .I1(inst92_O), .I2(inst29_O[7]), .I3(1'b0), .O(inst93_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst94 (.I0(inst2_Q), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst94_O));
SB_DFF inst95 (.C(CLKIN), .D(inst2_Q), .Q(inst95_Q));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst96 (.I0(inst2_Q), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst96_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst97 (.I0(inst95_Q), .I1(inst96_O), .I2(1'b0), .I3(1'b0), .O(inst97_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst98 (.I0(inst100_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst98_O));
Invert4 inst99 (.I({1'b1,1'b0,1'b0,1'b1}), .O(inst99_O));
Addcout4 inst100 (.I0(inst105_O), .I1(inst99_O), .O(inst100_O), .COUT(inst100_COUT));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst101 (.I0(inst102_O), .I1(inst97_O), .I2(1'b0), .I3(1'b0), .O(inst101_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst102 (.I0(inst98_O), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst102_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst103 (.I0(inst104_O), .I1(inst101_O), .I2(1'b0), .I3(1'b0), .O(inst103_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst104 (.I0(inst98_O), .I1(inst93_O), .I2(1'b0), .I3(1'b0), .O(inst104_O));
Counter4CER inst105 (.O(inst105_O), .COUT(inst105_COUT), .CLK(CLKIN), .CE(inst103_O), .RESET(inst108_O));
SB_LUT4 #(.LUT_INIT(16'h0400)) inst106 (.I0(inst105_O[0]), .I1(inst105_O[1]), .I2(inst105_O[2]), .I3(inst105_O[3]), .O(inst106_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst107 (.I0(inst106_O), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst107_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst108 (.I0(inst107_O), .I1(inst103_O), .I2(1'b0), .I3(1'b0), .O(inst108_O));
SIPO10CE inst109 (.I(inst2_Q), .O(inst109_O), .CLK(CLKIN), .CE(inst103_O));
SB_RAM40_4K #(.INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.READ_MODE(1),
.INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.WRITE_MODE(1),
.INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000)) inst110 (.RDATA(inst110_RDATA), .RADDR({1'b0,1'b0,inst25_O[8],inst25_O[7],inst25_O[6],inst25_O[5],inst25_O[4],inst25_O[3],inst25_O[2],inst25_O[1],inst25_O[0]}), .RCLK(CLKIN), .RCLKE(1'b1), .RE(1'b1), .WCLK(CLKIN), .WCLKE(1'b1), .WE(inst101_O), .WADDR({1'b0,1'b0,inst145_O[8],inst145_O[7],inst145_O[6],inst145_O[5],inst145_O[4],inst145_O[3],inst145_O[2],inst145_O[1],inst145_O[0]}), .MASK({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .WDATA({1'b0,inst109_O[8],1'b0,inst109_O[7],1'b0,inst109_O[6],1'b0,inst109_O[5],1'b0,inst109_O[4],1'b0,inst109_O[3],1'b0,inst109_O[2],1'b0,inst109_O[1]}));
Counter8CER inst111 (.O(inst111_O), .COUT(inst111_COUT), .CLK(CLKIN), .CE(inst101_O), .RESET(inst144_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst112 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst112_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst113 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst113_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst114 (.I0(inst112_O), .I1(inst113_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst114_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst115 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst115_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst116 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst116_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst117 (.I0(inst115_O), .I1(inst116_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst117_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst118 (.I0(inst114_O), .I1(inst117_O), .I2(inst111_O[5]), .I3(1'b0), .O(inst118_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst119 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst119_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst120 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst120_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst121 (.I0(inst119_O), .I1(inst120_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst121_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst122 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst122_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst123 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst123_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst124 (.I0(inst122_O), .I1(inst123_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst124_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst125 (.I0(inst121_O), .I1(inst124_O), .I2(inst111_O[5]), .I3(1'b0), .O(inst125_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst126 (.I0(inst118_O), .I1(inst125_O), .I2(inst111_O[6]), .I3(1'b0), .O(inst126_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst127 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst127_O));
SB_LUT4 #(.LUT_INIT(16'h0020)) inst128 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst128_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst129 (.I0(inst127_O), .I1(inst128_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst129_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst130 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst130_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst131 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst131_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst132 (.I0(inst130_O), .I1(inst131_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst132_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst133 (.I0(inst129_O), .I1(inst132_O), .I2(inst111_O[5]), .I3(1'b0), .O(inst133_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst134 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst134_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst135 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst135_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst136 (.I0(inst134_O), .I1(inst135_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst136_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst137 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst137_O));
SB_LUT4 #(.LUT_INIT(16'h0000)) inst138 (.I0(inst111_O[0]), .I1(inst111_O[1]), .I2(inst111_O[2]), .I3(inst111_O[3]), .O(inst138_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst139 (.I0(inst137_O), .I1(inst138_O), .I2(inst111_O[4]), .I3(1'b0), .O(inst139_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst140 (.I0(inst136_O), .I1(inst139_O), .I2(inst111_O[5]), .I3(1'b0), .O(inst140_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst141 (.I0(inst133_O), .I1(inst140_O), .I2(inst111_O[6]), .I3(1'b0), .O(inst141_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst142 (.I0(inst126_O), .I1(inst141_O), .I2(inst111_O[7]), .I3(1'b0), .O(inst142_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst143 (.I0(inst142_O), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst143_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst144 (.I0(inst143_O), .I1(inst101_O), .I2(1'b0), .I3(1'b0), .O(inst144_O));
Addcout9 inst145 (.I0({1'b0,inst111_O[7],inst111_O[6],inst111_O[5],inst111_O[4],inst111_O[3],inst111_O[2],inst111_O[1],inst111_O[0]}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .O(inst145_O), .COUT(inst145_COUT));
Mux2x4 inst146 (.I0({1'b0,1'b1,1'b0,1'b0}), .I1({1'b1,1'b0,1'b0,1'b1}), .S(inst16_O), .O(inst146_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst147 (.I0(inst149_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst147_O));
Invert4 inst148 (.I(inst146_O), .O(inst148_O));
Addcout4 inst149 (.I0(inst3_O), .I1(inst148_O), .O(inst149_O), .COUT(inst149_COUT));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst150 (.I0(inst147_O), .I1(inst10_Q), .I2(1'b0), .I3(1'b0), .O(inst150_O));
assign D4 = 1'b0;
assign D5 = 1'b0;
assign D6 = 1'b0;
assign D7 = 1'b0;
assign I = inst150_O;
assign D3 = 1'b0;
assign D2 = RX;
assign D1 = inst150_O;
assign D0 = inst2_Q;
endmodule

