module Addcout4 (input [3:0] I0, input [3:0] I1, output [3:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
assign O = {inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst7_CO;
endmodule

module Register4 (input [3:0] I, output [3:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
assign O = {inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter4 (output [3:0] O, output  COUT, input  CLK);
wire [3:0] inst0_O;
wire  inst0_COUT;
wire [3:0] inst1_O;
Addcout4 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register4 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout7 (input [6:0] I0, input [6:0] I1, output [6:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
assign O = {inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst13_CO;
endmodule

module Register7CE (input [6:0] I, output [6:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(I[6]), .Q(inst6_Q));
assign O = {inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter7CE (output [6:0] O, output  COUT, input  CLK, input  CE);
wire [6:0] inst0_O;
wire  inst0_COUT;
wire [6:0] inst1_O;
Addcout7 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register7CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Mux2x8 (input [7:0] I0, input [7:0] I1, input  S, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(S), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(S), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(S), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(S), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(I0[4]), .I1(I1[4]), .I2(S), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(I0[5]), .I1(I1[5]), .I2(S), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(I0[6]), .I1(I1[6]), .I2(S), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(I0[7]), .I1(I1[7]), .I2(S), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Addcout3 (input [2:0] I0, input [2:0] I1, output [2:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
assign O = {inst4_O,inst2_O,inst0_O};
assign COUT = inst5_CO;
endmodule

module Register3CE (input [2:0] I, output [2:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
assign O = {inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter3CE (output [2:0] O, output  COUT, input  CLK, input  CE);
wire [2:0] inst0_O;
wire  inst0_COUT;
wire [2:0] inst1_O;
Addcout3 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register3CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout8 (input [7:0] I0, input [7:0] I1, output [7:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
assign O = {inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst15_CO;
endmodule

module Register8CE (input [7:0] I, output [7:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter8CE (output [7:0] O, output  COUT, input  CLK, input  CE);
wire [7:0] inst0_O;
wire  inst0_COUT;
wire [7:0] inst1_O;
Addcout8 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register8CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Invert8 (input [7:0] I, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst4 (.I0(I[4]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst5 (.I0(I[5]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst6 (.I0(I[6]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(I[7]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Register3CER (input [2:0] I, output [2:0] O, input  CLK, input  CE, input  RESET);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
SB_DFFESR inst0 (.C(CLK), .R(RESET), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFESR inst1 (.C(CLK), .R(RESET), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFESR inst2 (.C(CLK), .R(RESET), .E(CE), .D(I[2]), .Q(inst2_Q));
assign O = {inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter3CER (output [2:0] O, output  COUT, input  CLK, input  CE, input  RESET);
wire [2:0] inst0_O;
wire  inst0_COUT;
wire [2:0] inst1_O;
Addcout3 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register3CER inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE), .RESET(RESET));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module PISO8CE (input  SI, input [7:0] PI, input  LOAD, output  O, input  CLK, input  CE);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire [7:0] inst8_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(SI), .I1(PI[0]), .I2(LOAD), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(inst8_O[0]), .I1(PI[1]), .I2(LOAD), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(inst8_O[1]), .I1(PI[2]), .I2(LOAD), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(inst8_O[2]), .I1(PI[3]), .I2(LOAD), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(inst8_O[3]), .I1(PI[4]), .I2(LOAD), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(inst8_O[4]), .I1(PI[5]), .I2(LOAD), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(inst8_O[5]), .I1(PI[6]), .I2(LOAD), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(inst8_O[6]), .I1(PI[7]), .I2(LOAD), .I3(1'b0), .O(inst7_O));
Register8CE inst8 (.I({inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O}), .O(inst8_O), .CLK(CLK), .CE(CE));
assign O = inst8_O[7];
endmodule

module Mux2x4 (input [3:0] I0, input [3:0] I1, input  S, output [3:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(S), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(S), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(S), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(S), .I3(1'b0), .O(inst3_O));
assign O = {inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Invert4 (input [3:0] I, output [3:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
assign O = {inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module main (output  I, output [4:0] J3, input  CLKIN);
wire [3:0] inst0_O;
wire  inst0_COUT;
wire [6:0] inst1_O;
wire  inst1_COUT;
wire [7:0] inst2_O;
wire [7:0] inst3_O;
wire [7:0] inst4_O;
wire [7:0] inst5_O;
wire [7:0] inst6_O;
wire [7:0] inst7_O;
wire [7:0] inst8_O;
wire [7:0] inst9_O;
wire [7:0] inst10_O;
wire [7:0] inst11_O;
wire [7:0] inst12_O;
wire [7:0] inst13_O;
wire [7:0] inst14_O;
wire [7:0] inst15_O;
wire [7:0] inst16_O;
wire [7:0] inst17_O;
wire [7:0] inst18_O;
wire [7:0] inst19_O;
wire [7:0] inst20_O;
wire [7:0] inst21_O;
wire [7:0] inst22_O;
wire [7:0] inst23_O;
wire [7:0] inst24_O;
wire [7:0] inst25_O;
wire [7:0] inst26_O;
wire [7:0] inst27_O;
wire [7:0] inst28_O;
wire [7:0] inst29_O;
wire [7:0] inst30_O;
wire [7:0] inst31_O;
wire [7:0] inst32_O;
wire [7:0] inst33_O;
wire [7:0] inst34_O;
wire [7:0] inst35_O;
wire [7:0] inst36_O;
wire [7:0] inst37_O;
wire [7:0] inst38_O;
wire [7:0] inst39_O;
wire [7:0] inst40_O;
wire [7:0] inst41_O;
wire [7:0] inst42_O;
wire [7:0] inst43_O;
wire [7:0] inst44_O;
wire [7:0] inst45_O;
wire [7:0] inst46_O;
wire [7:0] inst47_O;
wire [7:0] inst48_O;
wire [7:0] inst49_O;
wire [7:0] inst50_O;
wire [7:0] inst51_O;
wire [7:0] inst52_O;
wire [7:0] inst53_O;
wire [7:0] inst54_O;
wire [7:0] inst55_O;
wire [7:0] inst56_O;
wire [7:0] inst57_O;
wire [7:0] inst58_O;
wire [7:0] inst59_O;
wire [7:0] inst60_O;
wire [7:0] inst61_O;
wire [7:0] inst62_O;
wire [7:0] inst63_O;
wire [7:0] inst64_O;
wire [7:0] inst65_O;
wire [7:0] inst66_O;
wire [7:0] inst67_O;
wire [7:0] inst68_O;
wire [7:0] inst69_O;
wire [7:0] inst70_O;
wire [7:0] inst71_O;
wire [7:0] inst72_O;
wire [7:0] inst73_O;
wire [7:0] inst74_O;
wire [7:0] inst75_O;
wire [7:0] inst76_O;
wire [7:0] inst77_O;
wire [7:0] inst78_O;
wire [7:0] inst79_O;
wire [7:0] inst80_O;
wire [7:0] inst81_O;
wire [7:0] inst82_O;
wire [7:0] inst83_O;
wire [7:0] inst84_O;
wire [7:0] inst85_O;
wire [7:0] inst86_O;
wire [7:0] inst87_O;
wire [7:0] inst88_O;
wire [7:0] inst89_O;
wire [7:0] inst90_O;
wire [7:0] inst91_O;
wire [7:0] inst92_O;
wire [7:0] inst93_O;
wire [7:0] inst94_O;
wire [7:0] inst95_O;
wire [7:0] inst96_O;
wire [7:0] inst97_O;
wire [7:0] inst98_O;
wire [7:0] inst99_O;
wire [7:0] inst100_O;
wire [7:0] inst101_O;
wire [7:0] inst102_O;
wire [7:0] inst103_O;
wire [7:0] inst104_O;
wire [7:0] inst105_O;
wire [7:0] inst106_O;
wire [7:0] inst107_O;
wire [7:0] inst108_O;
wire [7:0] inst109_O;
wire [7:0] inst110_O;
wire [7:0] inst111_O;
wire [7:0] inst112_O;
wire [7:0] inst113_O;
wire [7:0] inst114_O;
wire [7:0] inst115_O;
wire [7:0] inst116_O;
wire [7:0] inst117_O;
wire [7:0] inst118_O;
wire [7:0] inst119_O;
wire [7:0] inst120_O;
wire [7:0] inst121_O;
wire [7:0] inst122_O;
wire [7:0] inst123_O;
wire [7:0] inst124_O;
wire [7:0] inst125_O;
wire [7:0] inst126_O;
wire [7:0] inst127_O;
wire [7:0] inst128_O;
wire [2:0] inst129_O;
wire  inst129_COUT;
wire  inst130_O;
wire [7:0] inst131_O;
wire  inst131_COUT;
wire  inst132_O;
wire [7:0] inst133_O;
wire [7:0] inst134_O;
wire  inst134_COUT;
wire  inst135_Q;
wire [2:0] inst136_O;
wire  inst136_COUT;
wire  inst137_O;
wire  inst138_Q;
wire  inst139_O;
wire  inst140_O;
wire  inst141_O;
wire  inst142_O;
wire  inst143_O;
wire [3:0] inst144_O;
wire  inst145_O;
wire [3:0] inst146_O;
wire [3:0] inst147_O;
wire  inst147_COUT;
wire  inst148_O;
Counter4 inst0 (.O(inst0_O), .COUT(inst0_COUT), .CLK(CLKIN));
Counter7CE inst1 (.O(inst1_O), .COUT(inst1_COUT), .CLK(CLKIN), .CE(inst143_O));
Mux2x8 inst2 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst2_O));
Mux2x8 inst3 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst3_O));
Mux2x8 inst4 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst4_O));
Mux2x8 inst5 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0}), .S(inst1_O[0]), .O(inst5_O));
Mux2x8 inst6 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst6_O));
Mux2x8 inst7 (.I0({1'b0,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst7_O));
Mux2x8 inst8 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1}), .S(inst1_O[0]), .O(inst8_O));
Mux2x8 inst9 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst9_O));
Mux2x8 inst10 (.I0({1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst10_O));
Mux2x8 inst11 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b0,1'b1,1'b1,1'b0,1'b1,1'b1}), .S(inst1_O[0]), .O(inst11_O));
Mux2x8 inst12 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst12_O));
Mux2x8 inst13 (.I0({1'b0,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst13_O));
Mux2x8 inst14 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0}), .S(inst1_O[0]), .O(inst14_O));
Mux2x8 inst15 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .S(inst1_O[0]), .O(inst15_O));
Mux2x8 inst16 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst16_O));
Mux2x8 inst17 (.I0({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst17_O));
Mux2x8 inst18 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .S(inst1_O[0]), .O(inst18_O));
Mux2x8 inst19 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst19_O));
Mux2x8 inst20 (.I0({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst20_O));
Mux2x8 inst21 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst21_O));
Mux2x8 inst22 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst22_O));
Mux2x8 inst23 (.I0({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst23_O));
Mux2x8 inst24 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .S(inst1_O[0]), .O(inst24_O));
Mux2x8 inst25 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst25_O));
Mux2x8 inst26 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst26_O));
Mux2x8 inst27 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst27_O));
Mux2x8 inst28 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst1_O[0]), .O(inst28_O));
Mux2x8 inst29 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst29_O));
Mux2x8 inst30 (.I0({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst30_O));
Mux2x8 inst31 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .S(inst1_O[0]), .O(inst31_O));
Mux2x8 inst32 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst32_O));
Mux2x8 inst33 (.I0({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst33_O));
Mux2x8 inst34 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst1_O[0]), .O(inst34_O));
Mux2x8 inst35 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst35_O));
Mux2x8 inst36 (.I0({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst36_O));
Mux2x8 inst37 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst37_O));
Mux2x8 inst38 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst38_O));
Mux2x8 inst39 (.I0({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst39_O));
Mux2x8 inst40 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst40_O));
Mux2x8 inst41 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst41_O));
Mux2x8 inst42 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst42_O));
Mux2x8 inst43 (.I0({1'b0,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst43_O));
Mux2x8 inst44 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1}), .S(inst1_O[0]), .O(inst44_O));
Mux2x8 inst45 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst45_O));
Mux2x8 inst46 (.I0({1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst46_O));
Mux2x8 inst47 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0}), .S(inst1_O[0]), .O(inst47_O));
Mux2x8 inst48 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst48_O));
Mux2x8 inst49 (.I0({1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst49_O));
Mux2x8 inst50 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0}), .S(inst1_O[0]), .O(inst50_O));
Mux2x8 inst51 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst51_O));
Mux2x8 inst52 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst52_O));
Mux2x8 inst53 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst53_O));
Mux2x8 inst54 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1}), .S(inst1_O[0]), .O(inst54_O));
Mux2x8 inst55 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst55_O));
Mux2x8 inst56 (.I0({1'b0,1'b0,1'b1,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst56_O));
Mux2x8 inst57 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst57_O));
Mux2x8 inst58 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst58_O));
Mux2x8 inst59 (.I0({1'b0,1'b1,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst59_O));
Mux2x8 inst60 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b0,1'b1,1'b0,1'b1,1'b1,1'b0}), .S(inst1_O[0]), .O(inst60_O));
Mux2x8 inst61 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst61_O));
Mux2x8 inst62 (.I0({1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst62_O));
Mux2x8 inst63 (.I0({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .I1({1'b0,1'b1,1'b1,1'b1,1'b0,1'b1,1'b0,1'b1}), .S(inst1_O[0]), .O(inst63_O));
Mux2x8 inst64 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .S(inst1_O[0]), .O(inst64_O));
Mux2x8 inst65 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst1_O[0]), .O(inst65_O));
Mux2x8 inst66 (.I0(inst2_O), .I1(inst3_O), .S(inst1_O[1]), .O(inst66_O));
Mux2x8 inst67 (.I0(inst4_O), .I1(inst5_O), .S(inst1_O[1]), .O(inst67_O));
Mux2x8 inst68 (.I0(inst6_O), .I1(inst7_O), .S(inst1_O[1]), .O(inst68_O));
Mux2x8 inst69 (.I0(inst8_O), .I1(inst9_O), .S(inst1_O[1]), .O(inst69_O));
Mux2x8 inst70 (.I0(inst10_O), .I1(inst11_O), .S(inst1_O[1]), .O(inst70_O));
Mux2x8 inst71 (.I0(inst12_O), .I1(inst13_O), .S(inst1_O[1]), .O(inst71_O));
Mux2x8 inst72 (.I0(inst14_O), .I1(inst15_O), .S(inst1_O[1]), .O(inst72_O));
Mux2x8 inst73 (.I0(inst16_O), .I1(inst17_O), .S(inst1_O[1]), .O(inst73_O));
Mux2x8 inst74 (.I0(inst18_O), .I1(inst19_O), .S(inst1_O[1]), .O(inst74_O));
Mux2x8 inst75 (.I0(inst20_O), .I1(inst21_O), .S(inst1_O[1]), .O(inst75_O));
Mux2x8 inst76 (.I0(inst22_O), .I1(inst23_O), .S(inst1_O[1]), .O(inst76_O));
Mux2x8 inst77 (.I0(inst24_O), .I1(inst25_O), .S(inst1_O[1]), .O(inst77_O));
Mux2x8 inst78 (.I0(inst26_O), .I1(inst27_O), .S(inst1_O[1]), .O(inst78_O));
Mux2x8 inst79 (.I0(inst28_O), .I1(inst29_O), .S(inst1_O[1]), .O(inst79_O));
Mux2x8 inst80 (.I0(inst30_O), .I1(inst31_O), .S(inst1_O[1]), .O(inst80_O));
Mux2x8 inst81 (.I0(inst32_O), .I1(inst33_O), .S(inst1_O[1]), .O(inst81_O));
Mux2x8 inst82 (.I0(inst34_O), .I1(inst35_O), .S(inst1_O[1]), .O(inst82_O));
Mux2x8 inst83 (.I0(inst36_O), .I1(inst37_O), .S(inst1_O[1]), .O(inst83_O));
Mux2x8 inst84 (.I0(inst38_O), .I1(inst39_O), .S(inst1_O[1]), .O(inst84_O));
Mux2x8 inst85 (.I0(inst40_O), .I1(inst41_O), .S(inst1_O[1]), .O(inst85_O));
Mux2x8 inst86 (.I0(inst42_O), .I1(inst43_O), .S(inst1_O[1]), .O(inst86_O));
Mux2x8 inst87 (.I0(inst44_O), .I1(inst45_O), .S(inst1_O[1]), .O(inst87_O));
Mux2x8 inst88 (.I0(inst46_O), .I1(inst47_O), .S(inst1_O[1]), .O(inst88_O));
Mux2x8 inst89 (.I0(inst48_O), .I1(inst49_O), .S(inst1_O[1]), .O(inst89_O));
Mux2x8 inst90 (.I0(inst50_O), .I1(inst51_O), .S(inst1_O[1]), .O(inst90_O));
Mux2x8 inst91 (.I0(inst52_O), .I1(inst53_O), .S(inst1_O[1]), .O(inst91_O));
Mux2x8 inst92 (.I0(inst54_O), .I1(inst55_O), .S(inst1_O[1]), .O(inst92_O));
Mux2x8 inst93 (.I0(inst56_O), .I1(inst57_O), .S(inst1_O[1]), .O(inst93_O));
Mux2x8 inst94 (.I0(inst58_O), .I1(inst59_O), .S(inst1_O[1]), .O(inst94_O));
Mux2x8 inst95 (.I0(inst60_O), .I1(inst61_O), .S(inst1_O[1]), .O(inst95_O));
Mux2x8 inst96 (.I0(inst62_O), .I1(inst63_O), .S(inst1_O[1]), .O(inst96_O));
Mux2x8 inst97 (.I0(inst64_O), .I1(inst65_O), .S(inst1_O[1]), .O(inst97_O));
Mux2x8 inst98 (.I0(inst66_O), .I1(inst67_O), .S(inst1_O[2]), .O(inst98_O));
Mux2x8 inst99 (.I0(inst68_O), .I1(inst69_O), .S(inst1_O[2]), .O(inst99_O));
Mux2x8 inst100 (.I0(inst70_O), .I1(inst71_O), .S(inst1_O[2]), .O(inst100_O));
Mux2x8 inst101 (.I0(inst72_O), .I1(inst73_O), .S(inst1_O[2]), .O(inst101_O));
Mux2x8 inst102 (.I0(inst74_O), .I1(inst75_O), .S(inst1_O[2]), .O(inst102_O));
Mux2x8 inst103 (.I0(inst76_O), .I1(inst77_O), .S(inst1_O[2]), .O(inst103_O));
Mux2x8 inst104 (.I0(inst78_O), .I1(inst79_O), .S(inst1_O[2]), .O(inst104_O));
Mux2x8 inst105 (.I0(inst80_O), .I1(inst81_O), .S(inst1_O[2]), .O(inst105_O));
Mux2x8 inst106 (.I0(inst82_O), .I1(inst83_O), .S(inst1_O[2]), .O(inst106_O));
Mux2x8 inst107 (.I0(inst84_O), .I1(inst85_O), .S(inst1_O[2]), .O(inst107_O));
Mux2x8 inst108 (.I0(inst86_O), .I1(inst87_O), .S(inst1_O[2]), .O(inst108_O));
Mux2x8 inst109 (.I0(inst88_O), .I1(inst89_O), .S(inst1_O[2]), .O(inst109_O));
Mux2x8 inst110 (.I0(inst90_O), .I1(inst91_O), .S(inst1_O[2]), .O(inst110_O));
Mux2x8 inst111 (.I0(inst92_O), .I1(inst93_O), .S(inst1_O[2]), .O(inst111_O));
Mux2x8 inst112 (.I0(inst94_O), .I1(inst95_O), .S(inst1_O[2]), .O(inst112_O));
Mux2x8 inst113 (.I0(inst96_O), .I1(inst97_O), .S(inst1_O[2]), .O(inst113_O));
Mux2x8 inst114 (.I0(inst98_O), .I1(inst99_O), .S(inst1_O[3]), .O(inst114_O));
Mux2x8 inst115 (.I0(inst100_O), .I1(inst101_O), .S(inst1_O[3]), .O(inst115_O));
Mux2x8 inst116 (.I0(inst102_O), .I1(inst103_O), .S(inst1_O[3]), .O(inst116_O));
Mux2x8 inst117 (.I0(inst104_O), .I1(inst105_O), .S(inst1_O[3]), .O(inst117_O));
Mux2x8 inst118 (.I0(inst106_O), .I1(inst107_O), .S(inst1_O[3]), .O(inst118_O));
Mux2x8 inst119 (.I0(inst108_O), .I1(inst109_O), .S(inst1_O[3]), .O(inst119_O));
Mux2x8 inst120 (.I0(inst110_O), .I1(inst111_O), .S(inst1_O[3]), .O(inst120_O));
Mux2x8 inst121 (.I0(inst112_O), .I1(inst113_O), .S(inst1_O[3]), .O(inst121_O));
Mux2x8 inst122 (.I0(inst114_O), .I1(inst115_O), .S(inst1_O[4]), .O(inst122_O));
Mux2x8 inst123 (.I0(inst116_O), .I1(inst117_O), .S(inst1_O[4]), .O(inst123_O));
Mux2x8 inst124 (.I0(inst118_O), .I1(inst119_O), .S(inst1_O[4]), .O(inst124_O));
Mux2x8 inst125 (.I0(inst120_O), .I1(inst121_O), .S(inst1_O[4]), .O(inst125_O));
Mux2x8 inst126 (.I0(inst122_O), .I1(inst123_O), .S(inst1_O[5]), .O(inst126_O));
Mux2x8 inst127 (.I0(inst124_O), .I1(inst125_O), .S(inst1_O[5]), .O(inst127_O));
Mux2x8 inst128 (.I0(inst126_O), .I1(inst127_O), .S(inst1_O[6]), .O(inst128_O));
Counter3CE inst129 (.O(inst129_O), .COUT(inst129_COUT), .CLK(CLKIN), .CE(inst0_COUT));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst130 (.I0(inst0_COUT), .I1(inst129_COUT), .I2(1'b0), .I3(1'b0), .O(inst130_O));
Counter8CE inst131 (.O(inst131_O), .COUT(inst131_COUT), .CLK(CLKIN), .CE(inst130_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst132 (.I0(inst134_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst132_O));
Invert8 inst133 (.I({1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}), .O(inst133_O));
Addcout8 inst134 (.I0(inst131_O), .I1(inst133_O), .O(inst134_O), .COUT(inst134_COUT));
SB_DFFE inst135 (.C(CLKIN), .E(inst0_COUT), .D(inst132_O), .Q(inst135_Q));
Counter3CER inst136 (.O(inst136_O), .COUT(inst136_COUT), .CLK(CLKIN), .CE(inst0_COUT), .RESET(inst140_O));
SB_LUT4 #(.LUT_INIT(16'h0080)) inst137 (.I0(inst136_O[0]), .I1(inst136_O[1]), .I2(inst136_O[2]), .I3(1'b0), .O(inst137_O));
SB_DFFE inst138 (.C(CLKIN), .E(inst0_COUT), .D(inst139_O), .Q(inst138_Q));
SB_LUT4 #(.LUT_INIT(16'h5454)) inst139 (.I0(inst137_O), .I1(inst132_O), .I2(inst138_Q), .I3(1'b0), .O(inst139_O));
SB_LUT4 #(.LUT_INIT(16'h2222)) inst140 (.I0(inst137_O), .I1(inst138_Q), .I2(1'b0), .I3(1'b0), .O(inst140_O));
PISO8CE inst141 (.SI(1'b1), .PI(inst128_O), .LOAD(inst142_O), .O(inst141_O), .CLK(CLKIN), .CE(inst0_COUT));
SB_LUT4 #(.LUT_INIT(16'h2222)) inst142 (.I0(inst132_O), .I1(inst138_Q), .I2(1'b0), .I3(1'b0), .O(inst142_O));
SB_LUT4 #(.LUT_INIT(16'h4444)) inst143 (.I0(inst138_Q), .I1(inst0_COUT), .I2(1'b0), .I3(1'b0), .O(inst143_O));
Mux2x4 inst144 (.I0({1'b0,1'b1,1'b0,1'b0}), .I1({1'b1,1'b0,1'b0,1'b1}), .S(inst141_O), .O(inst144_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst145 (.I0(inst147_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst145_O));
Invert4 inst146 (.I(inst144_O), .O(inst146_O));
Addcout4 inst147 (.I0(inst0_O), .I1(inst146_O), .O(inst147_O), .COUT(inst147_COUT));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst148 (.I0(inst145_O), .I1(inst135_Q), .I2(1'b0), .I3(1'b0), .O(inst148_O));
assign I = inst148_O;
assign J3 = {inst148_O,inst138_Q,inst135_Q,inst0_COUT,1'b0};
endmodule

